// modulo transmissor UART

module tx(
    input  logic clk,        
    input  logic tick,       // Tick de baud rate (ex: 9600Hz)
    input  logic send,       // Sinal para iniciar transmissão
    input  logic [7:0]  data_in, // Byte de dados
    output logic tx,         // Linha TX
    output logic busy        // Indica transmissão em andamento
);

    logic [3:0] bit_cnt = 0;
    logic [9:0] shift_reg = 10'b1111111111;  // Linha ociosa = 1
    logic sending = 0;

    // Função para calcular paridade par
    function logic calc_parity(input [7:0] data);
        calc_parity = ~^data;  // XOR de todos os bits e inverte (paridade par)
    endfunction

    always_ff @(posedge clk) begin
        if (send && !sending) begin
            shift_reg <= {1'b1,  data_in,  calc_parity(data_in), 1'b0}; // STOP | PAR | DATA | START
            bit_cnt   <= 0;
            sending   <= 1;
            busy      <= 1;
            tx        <= 0; // START bit
        end
        else if (tick && sending) begin
            tx        <= shift_reg[0];
            shift_reg <= shift_reg >> 1;
            bit_cnt   <= bit_cnt + 1;

            if (bit_cnt == 9) begin
                sending <= 0;
                busy    <= 0;
                tx      <= 1; // Linha idle após fim
            end
        end else if (!sending) begin
            tx <= 1; // idle
        end
    end


endmodule