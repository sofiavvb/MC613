// clock para board -> unit watch e stopwatch

module clock (
    input logic CLOCK_50,
    input logic[3:0] KEY,


);








endmodule
